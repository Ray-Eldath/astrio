package ALUType;
    typedef enum bit [3:0]{
        AND, OR, ADD, SUB, LESS_THAN, XOR
    } cmd_t /* verilator public */;
endpackage : ALUType