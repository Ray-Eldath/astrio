package Types;
    typedef logic unsigned [31:0] addr_t;

    typedef logic signed [31:0] op_t;
    typedef reg signed [31:0] op_reg_t;
    typedef logic unsigned [4:0] reg_id_t;

    typedef logic unsigned [31:0] inst_t;
    typedef reg unsigned [31:0] inst_reg_t;
endpackage : Types