package Parameters;
    parameter InstSpace/* verilator public */=1024;
    parameter InstStartFrom /* verilator public */=32'h0040_0000;
endpackage : Parameters
