package PCType;
    typedef enum bit [1:0]{
        NONE, INC, LOAD
    } cmd_t /* verilator public */;
endpackage : PCType