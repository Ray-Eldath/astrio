package Types;
    typedef bit unsigned [31:0] addr_t;

    typedef bit signed [31:0] op_t;
    typedef bit unsigned [4:0] reg_id_t;

    typedef bit unsigned [31:0] inst_t;
endpackage : Types