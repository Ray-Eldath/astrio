package Mux3Type;
    typedef enum bit [1:0]{
        ZERO, DEFAULT, LEFT, RIGHT
    } cmd_t;
endpackage : Mux3Type