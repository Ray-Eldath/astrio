package PCType;
    typedef enum bit [1:0]{
        NONE, INC, LOAD
    } pc_cmd_t /* verilator public */;
endpackage : PCType