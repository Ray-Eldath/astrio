package Mux3Type;
    typedef enum bit [1:0]{
        DEFAULT, TOP, BOTTOM, ZERO
    } cmd_t;
endpackage : Mux3Type